package tta0_params is
  constant fu_LSU_dataw : integer := 32;
  constant fu_LSU_addrw : integer := 24;
  constant fu_INPUT_statusw : integer := 9;
  constant fu_OUTPUT_statusw : integer := 9;
end tta0_params;
